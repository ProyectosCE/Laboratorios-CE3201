module ALU_N_bits 
	#(parameter N=4)
	 (input logic[N-1:0] a, b,
	  input logic[1:0] control, // 2 bits for 4 op, need 
	  output logic[N-1:0] result,
	  output logic v, c, n, z);
	// Wires
	
	// Operations
		// OR
		// AND
		// Add
		1. codigo
			- maquina (ALU)
			- operaciones
				and 
				or 
				- 
				+ 
				
				*
				/
				%
				<<
				>>
				xor
				
				xor
		
		
		2. timming
			- Leer
			
		
		// Sub
		or()
		and()
		xor(a,b)
	// Mux
	
	// Flags
	



endmodule
